library verilog;
use verilog.vl_types.all;
entity gpul_vlg_vec_tst is
end gpul_vlg_vec_tst;
